* Definindo a temperatura de operação
.TEMP 25

* Declarando parametros que serão utilizados nas simulações

.include 32LP.mod
.include 32HP.mod

* Declarando parametros que serão utilizados nas simulações
.param supply = 0.9

* Declaração das fontes
vdd source 0 dc 0.9
venable enable 0 PWL(0 0.9) r=-1
*vclock 7 5 PWL(0 1 20ns 0) r=-1

* NAND 
MP1 out_nand enable        source   source PMOS_32HP L=32n W=100n
MP2 out_nand out_oscilador source   source PMOS_32HP L=32n W=100n
MN1 out_nand enable        dnmos    0      NMOS_32HP L=32n W=100n
MN2 dnmos    out_oscilador 0        0      NMOS_32HP L=32n W=100n  


* Declaração do inversor 1
MP_hp1 out_inv1 out_nand source source PMOS_32HP L=32n W=100n
MN_hp1 out_inv1 out_nand 0      0      NMOS_32HP L=32n W=100n

* Declaração do inversor 2
MP_hp2 out_inv2 out_inv1 source source PMOS_32HP L=32n W=100n
MN_hp2 out_inv2 out_inv1 0      0      NMOS_32HP L=32n W=100n

* Declaração do inversor 3
MP_hp3 out_inv3 out_inv2 source source PMOS_32HP L=32n W=100n
MN_hp3 out_inv3 out_inv2 0      0      NMOS_32HP L=32n W=100n

* Declaração do inversor 4
MP_hp4 out_inv4 out_inv3 source source PMOS_32HP L=32n W=100n
MN_hp4 out_inv4 out_inv3 0      0      NMOS_32HP L=32n W=100n

* Declaração do inversor 5
MP_hp5 out_inv5 out_inv4 source source PMOS_32HP L=32n W=100n
MN_hp5 out_inv5 out_inv4 0      0      NMOS_32HP L=32n W=100n

* Declaração do inversor 6
MP_hp6 out_inv6 out_inv5 source source PMOS_32HP L=32n W=100n
MN_hp6 out_inv6 out_inv5 0      0      NMOS_32HP L=32n W=100n

* Declaração do inversor 7
MP_hp7 out_inv7 out_inv6 source source PMOS_32HP L=32n W=100n
MN_hp7 out_inv7 out_inv6 0      0      NMOS_32HP L=32n W=100n

* Declaração do inversor 8
MP_hp8 out_inv8 out_inv7 source source PMOS_32HP L=32n W=100n
MN_hp8 out_inv8 out_inv7 0      0      NMOS_32HP L=32n W=100n
* Declaração do inversor 9
MP_hp9 out_inv9 out_inv8 source source PMOS_32HP L=32n W=100n
MN_hp9 out_inv9 out_inv8 0      0      NMOS_32HP L=32n W=100n
* Declaração do inversor 10
MP_hp10 out_inv10 out_inv9 source source PMOS_32HP L=32n W=100n
MN_hp10 out_inv10 out_inv9 0      0      NMOS_32HP L=32n W=100n
* Declaração do inversor 11
MP_hp11 out_inv11 out_inv10 source source PMOS_32HP L=32n W=100n
MN_hp11 out_inv11 out_inv10 0      0      NMOS_32HP L=32n W=100n
* Declaração do inversor 12
MP_hp12 out_inv12 out_inv11 source source PMOS_32HP L=32n W=100n
MN_hp12 out_inv12 out_inv11 0      0      NMOS_32HP L=32n W=100n
* Declaração do inversor 13
MP_hp13 out_inv13 out_inv12 source source PMOS_32HP L=32n W=100n
MN_hp13 out_inv13 out_inv12 0      0      NMOS_32HP L=32n W=100n
* Declaração do inversor 14
MP_hp14 out_inv14 out_inv13 source source PMOS_32HP L=32n W=100n
MN_hp14 out_inv14 out_inv13 0      0      NMOS_32HP L=32n W=100n
* Declaração do inversor 15
MP_hp15 out_inv15 out_inv14 source source PMOS_32HP L=32n W=100n
MN_hp15 out_inv15 out_inv14 0      0      NMOS_32HP L=32n W=100n
* Declaração do inversor 16
MP_hp16 out_oscilador out_inv15 source source PMOS_32HP L=32n W=100n
MN_hp16 out_oscilador out_inv15 0      0      NMOS_32HP L=32n W=100n


* Declarando o tipo de simulação 

.tran 0.005n 1n
*******************************************************************

.control

run

* saida lógica
*spec 0 1K 100 3

    set color0=white
    set xbrushwidth=3

    plot v(out_oscilador) 
    plot v(out_oscilador) v(enable)
    
.endc
.end