* Definindo a temperatura de operação
.TEMP 25

* Declarando parametros que serão utilizados nas simulações

.include 32HP.mod

* Declarando parametros que serão utilizados nas simulações
.param supply = 0.9

* Declaração das fontes
vdd vdd 0 dc 1.8
vin1 in1 0 PULSE (0 1.8 0 0.1n 0.1n 5n 10n)
vin2 in2 0 PULSE (0 1.8 0 0.1n 0.1n 10n 20n)





* NAND 

MP1 out in1 vpmos vdd PMOS_32HP L=32n W=100n
MP2 out in2 vpmos vdd PMOS_32HP L=32n W=100n
MN1 out in1 dnmos 0 NMOS_32HP L=32n W=100n
MN2 dnmos in2 0 0 NMOS_32HP L=32n W=100n


* Declarando o tipo de simulação 

* Declarando o tipo de simulação 
.dc vinput 0 0.9 0.01

.control

run

* saida lógica
*spec 0 1K 100 3

    set color0=white
    set xbrushwidth=3

    plot v(in1)
    plot v(in2)
    plot v(in1) v(in2)
    plot i(vnmos) i(vpmos)

.endc
.end