* Simulação de um inversor
* Incluindo o modelo do Transistor 
.include 32HP.mod
.include 32LP.mod

* Definindo a temperatura de operação
.TEMP 25

* Declarando parametros que serão utilizados nas simulações
.param supply = 0.9

* Declaração das fontes
valimentacao vdd 0 supply
vinput in 0 0.45
vout out 0 0

vpmos dpmos out 0
vnmos out dnmos 0

vpmos_a out dpmos_a 0
vnmos_a out dnmos_a 0

* Declaração do inversor 32 high power
MP_hp vdd in out_32hp vdd PMOS_32HP L=32n W=200n
MN_hp 0   in out_32hp 0   NMOS_32HP L=32n W=100n

* Declaração do inversor 32 low peformance
MP_lp vdd in out_32lp vdd PMOS_32lp L=32n W=200n
MN_lp 0   in out_32lp 0   NMOS_32lp L=32n W=100n

* MPb vdd in dpmos vdd PMOS_32lp L=32n W=200n 
* MNb 0   in dnmos 0  NMOS_32lp L=32n W=100n

* Pa vdd in dpmos_a vdd PMOS_lp L=32n W=200n
* MNa 0   in dnmos_a 0   NMOS_lp L=32n W=100n

* Declarando o tipo de simulação 
* .DC <fonte_que_sofrerá_variação> <valor_inicial_da_variação> <valor_final_da_variação> <passo_da_variação>
.dc vinput 0 0.9 0.01
*.dc vout 0 0.9 0.01 vinput 0 0.9 0.15

*******************************************************************
* parametros de simulação

.control

run

* saidas lógicas
plot out_32hp out_32lp


.endc