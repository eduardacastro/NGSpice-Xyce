* Definindo a temperatura de operação
.TEMP 25

* Declarando parametros que serão utilizados nas simulações

.include 32LP.mod
.include 32HP.mod

* Declarando parametros que serão utilizados nas simulações
.param supply = 0.9

* Declaração das fontes
venable enable 0 PULSE (0 1.8 0 0.1n 0.1n 5n 10n)


* NAND 

MP1 out_nand enable vpmos vdd PMOS_32HP L=32n W=100n
MP2 out_nand out_oscilador vpmos vdd PMOS_32HP L=32n W=100n
MN1 out_nand enable dnmos 0 NMOS_32HP L=32n W=100n
MN2 dnmos out_oscilador 0 0 NMOS_32HP L=32n W=100n


* Declaração do inversor 1
MP_hp1 vdd out_nand out_inv1 vdd PMOS_32HP L=32n W=100n
MN_hp1 0   out_nand out_inv1 0   NMOS_32HP L=32n W=100n

* Declaração do inversor 2
MP_hp2 vdd out_inv1 out_inv2 vdd PMOS_32HP L=32n W=100n
MN_hp2 0   out_inv1 out_inv2 0   NMOS_32HP L=32n W=100n

* Declaração do inversor 3
MP_hp3 vdd out_inv2 out_inv3 vdd PMOS_32HP L=32n W=100n
MN_hp3 0   out_inv2 out_inv3 0   NMOS_32HP L=32n W=100n

* Declaração do inversor 4
MP_hp4 vdd out_inv3 out_oscilador vdd PMOS_32HP L=32n W=100n
MN_hp4 0   out_inv3 out_oscilador 0   NMOS_32HP L=32n W=100n


* Declarando o tipo de simulação 

.tran 0.1n 50n
*******************************************************************

.control

run

* saida lógica
*spec 0 1K 100 3

    set color0=white
    set xbrushwidth=3

    plot v(out_oscilador) 
    plot v(out_oscilador) v(enable)
    
.endc
.end