* Definindo a temperatura de operação
.TEMP 25

* Declarando parametros que serão utilizados nas simulações

.include 32LP.mod
.include 32HP.mod

* Declarando parametros que serão utilizados nas simulações
.param supply = 0.9

* Declaração das fontes
valimentacao vdd 0 supply
vinput in 0 0.45
vout out 0 0


* NAND 
** Paralelo
MP1 out_hp in vdd vdd PMOS_32HP L=32n W=100n
MP2 out_hp in vdd vdd PMOS_32HP L=32n W=100n
** Serie
MN1 out_hp in dnmos 0 NMOS_32HP L=32n W=100n
MN2 dnmos in 0 0 NMOS_32HP L=32n W=100n


MP1lp out_lp in vdd vdd PMOS_32LP L=32n W=100n
MP2lp out_lp in vdd vdd PMOS_32LP L=32n W=100n
** Serie
MN1lp out_lp in dnmos 0 NMOS_32LP L=32n W=100n
MN2lp dnmos in 0 0 NMOS_32LP L=32n W=100n


* Declarando o tipo de simulação 
.dc vinput 0 0.9 0.01
*******************************************************************
* parametros de simulação

.op
