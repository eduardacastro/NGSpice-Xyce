*  cd ../../Users/Asus/Desktop/NGSpice/ckt-inversor/Xyce
* Definindo a temperatura de operação
.param agingp = -0.16
.param agingn = 0.16
.include "finfet.mod"
.param supply = 0.7

* Declaração das fontes
vdd vdd 0 dc 0.7
vin1 in 0 PULSE (0 0.7 100p 10p 10p 100p 300p)
Vagingp1 inp1 in dc 0
Vagingn1 in inn1 dc 0
.tran 0.001p 1000p

 
MP1 out inp1 vdd vdd pmos_lvt L=20n NFIN=4
MN1 out inn1 0 0 nmos_lvt L=20n NFIN=4

cload out 0 0.5f

*vaux out aux 0
* Positivo
*iexp 0 aux exp(0 145u 150p 2p 165p 4p)
* Negativo
*iexp2 aux 0 exp(0 155u 550p 2p 565p 4p)

.PRINT TRAN FORMAT=CSV v(out) v(in)
.MEASURE TRAN HL TRIG v(in) VAL='supply*0.5' RISE=1 TARG v(out) VAL='supply*0.5' FALL=1 
.MEASURE TRAN LH TRIG v(in) VAL='supply*0.5' FALL=1 TARG v(out) VAL='supply*0.5' RISE=1 
.MEASURE TRAN Fall TRIG v(out) VAL='supply*0.8' FALL=1 TARG v(out) VAL='supply*0.2' FALL=1
.MEASURE TRAN RISE TRIG v(out) VAL='supply*0.2' RISE=1 TARG v(out) VAL='supply*0.8' RISE=1

*meas tran tp_hl_in1 trig v(in1) val=0.45 rise=1 targ v(out) val=0.45 fall=1
*meas tran tp_lh_in1 trig v(in1) val=0.45 fall=1 targ v(out) val=0.45 rise=1
*meas tran tp_fall_in1 trig v(out) val=0.72 fall=1 targ v(out) val=0.18 fall=1
*meas tran tp_rise_in1 trig v(out) val=0.18 rise=1 targ v(out) val=0.72 rise=1

.end