*  cd ../../NGSpice/ckt-aoi
* Definindo a temperatura de operação
.TEMP 25

* Declarando parametros que serão utilizados nas simulações
.param agingp = -0.01
.param agingn = 0.01
.param Wn = 100n
.param Wp = 200n
.param WnInv = 100n
.param WpInv = 200n
.include 32HP.mod
* Declaração das fontes
vdd vdd 0 dc 0.9

* Variando Inv1
*vin1 in1 0 PULSE (0 0.9 0p 10p 10p 300p 600p)
*vin2 in2 0 PULSE (0 0 0p 10p 10p 300p 600p)
*vin3 in3 0 PULSE (0 0 0p 10p 10p 300p 600p)

*Variando In2 e In3 usar esses 
vin1 in1 0 PULSE (0 0 300p 10p 10p 300p 600p)
vin3 in3 0 PULSE (0 0.9 0p 10p 10p 300p 600p)
vin2 in2 0 PULSE (0 0.9 0p 10p 10p 1200p 1200p)


Vagingp1 in1 inp1 dc agingp
Vagingn1 in1 inn1 dc agingn
Vagingp2 in2 inp2 dc agingp
Vagingn2 in2 inn2 dc agingn
Vagingp3 in3 inp3 dc agingp
Vagingn3 in3 inn3 dc agingn


MP1 saida inp1 vdd vdd PMOS_32HP L=32n W=Wp
MP3 out inp3 saida saida PMOS_32HP L=32n W=Wp
MP2 out inp2 saida saida PMOS_32HP L=32n W=Wp


MN1 out inn1 0 0 NMOS_32HP L=32n W=Wn
MN2 out inn2 dnmos dnmos NMOS_32HP L=32n W=Wn
MN3 dnmos inn3 0 0 NMOS_32HP L=32n W=Wn

*LOAD INV (FoF - Fanout of Four - emula 4 Invs usando sizing)
MPload outload out vdd vdd PMOS_32HP L=32n W=WpInv
MNload outload out 0 0 NMOS_32HP L=32n W=WnInv

MPloade1 outload1 outload vdd vdd PMOS_32HP L=32n W=WpInv
MNloade1 outload1 outload 0 0 NMOS_32HP L=32n W=WnInv

MPloade2 outload2 outload1 vdd vdd PMOS_32HP L=32n W=WpInv
MNloade2 outload2 outload1 0 0 NMOS_32HP L=32n W=WnInv

vaux out aux 0
* sinal positivo
iexp 0 aux exp(0 90u 750p 2p 765p 4p)
*sinal negativo0
iexp2 aux 0 exp(0 90u 450p 2p 465p 4p)
* Declarando o tipo de simulação 


*.tran 0.1p 500p
.tran 0.1p 900p
***********************
* parametros de simulação

.control

run
  set color0=gray
  set xbrushwidth=3
plot v(outload2)-3 v(outload1)-2 v(outload)-1 v(out) v(in1)+1 v(in2)+2 v(in3)+3 
*plot i(vaux)
*Variando Inv2
meas tran tp_hl_in2_in1_0 trig v(in3) val=0.45 rise=2 targ v(out) val=0.45 fall=2
meas tran tp_lh_in2_in1_0 trig v(in3) val=0.45 fall=1 targ v(out) val=0.45 rise=1
meas tran tp_fall_in2_in1_0 trig v(out) val=0.72 fall=2 targ v(out) val=0.18 fall=2
meas tran tp_rise_in2_in1_0 trig v(out) val=0.18 rise=1 targ v(out) val=0.72 rise=1

*Variando Inv1
*plot v(out) v(in1)+1 v(in2)+2 v(in3)+3 
*meas tran tp_hl_in1_in2_0 trig v(in1) val=0.45 rise=2 targ v(out) val=0.45 fall=2
*meas tran tp_lh_in1_in2_0 trig v(in1) val=0.45 fall=1 targ v(out) val=0.45 rise=1
*meas tran tp_fall_in1_in2_0 trig v(out) val=0.72 fall=2 targ v(out) val=0.18 fall=2
*meas tran tp_rise_in1_in2_0 trig v(out) val=0.18 rise=1 targ v(out) val=0.72 rise=1


.endc
.end