*  cd ../../Users/Asus/Desktop/NGSpice/ckt-nor/Xyce/nor-2
.include "finfet.mod"
* Declaração das fontes
.param supply = 0.7
vdd vdd 0 dc 0.7
vin1 in2 0 PULSE (0 0.0 100p 10p 10p 1000p 1000p)
vin2 in1 0 PULSE (0 0.7 0p 10p 10p 300p 500p)
vin3 in3 0 PULSE (0 0.0 100p 10p 10p 1000p 1000p)
.tran 0.001p 1000p
Vagingp1 in1 inp1 dc -0.0445
Vagingp2 in2 inp2 dc -0.0397
Vagingp3 in3 inp3 dc -0.0354
Vagingn1 in1 inn1 dc 0.0445
Vagingn2 in2 inn2 dc 0.0445
Vagingn3 in3 inn3 dc 0.0445


MP1 vpmos inp1 vdd vdd pmos_lvt L=20n NFIN=2
MP2 vp2mos inp2 vpmos vdd pmos_lvt L=20n NFIN=2 
MP3 out inp3 vp2mos vdd pmos_lvt L=20n NFIN=2 
MN1 out inn1 0 0 nmos_lvt L=20n NFIN=2 
MN2 out inn2 0 0 nmos_lvt L=20n NFIN=2
MN3 out inn3 0 0 nmos_lvt L=20n NFIN=2 

.OPTION OUTPUT INITIAL_INTERVAL=.1ps 350ps
.PRINT TRAN FORMAT=CSV v(out) v(in1) v(in2) v(in3)
*Variando Inv1
.MEASURE TRAN HL1 TRIG v(in1) VAL='supply*0.5' RISE=2 TARG v(out) VAL='supply*0.5' FALL=2
.MEASURE TRAN LH1 TRIG v(in1) VAL='supply*0.5' FALL=1 TARG v(out) VAL='supply*0.5' RISE=1

*Variando Inv2
.MEASURE TRAN HL2 TRIG v(in2) VAL='supply*0.5' RISE=2 TARG v(out) VAL='supply*0.5' FALL=2
.MEASURE TRAN LH2 TRIG v(in2) VAL='supply*0.5' FALL=1 TARG v(out) VAL='supply*0.5' RISE=1

*Variando Inv2
.MEASURE TRAN HL3 TRIG v(in3) VAL='supply*0.5' RISE=2 TARG v(out) VAL='supply*0.5' FALL=2
.MEASURE TRAN LH3 TRIG v(in3) VAL='supply*0.5' FALL=1 TARG v(out) VAL='supply*0.5' RISE=1 

.MEASURE TRAN Fall TRIG v(out) VAL='supply*0.8' FALL=2 TARG v(out) VAL='supply*0.2' FALL=2
.MEASURE TRAN RISE TRIG v(out) VAL='supply*0.2' RISE=2 TARG v(out) VAL='supply*0.8' RISE=2

.end