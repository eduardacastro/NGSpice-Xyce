*  cd ../../Users/Asus/Desktop/NGSpice/ckt-inversor/Xyce
* Definindo a temperatura de operação
.include "finfet.mod"
.param supply = 0.7

* Declaração das fontes
vdd vdd 0 dc 0.7
vin1 in 0 PULSE (0 0.7 100p 10p 10p 300p 600p)
Vagingp1 in inp1 dc -0.0445
Vagingn1 in inn1 dc 0.0445
.tran 0.001p 1000p

 
MP1 out in vdd vdd pmos_lvt L=20n NFIN=2
MN1 out in 0 0 nmos_lvt L=20n NFIN=2


vaux out aux 0
* Positivo
iexp 0 aux exp(0 65u 120p 2p 135p 4p)
* Negativo
iexp2 aux 0 exp(0 50u 440p 2p 455p 4p)


.OPTION OUTPUT INITIAL_INTERVAL=.01ps 0.350ps
.PRINT TRAN FORMAT=CSV v(out) v(in)

.end