* Definindo a temperatura de operação
.TEMP 25

* Declarando parametros que serão utilizados nas simulações


.include 32HP.mod

* Declaração das fontes
vdd vdd 0 0v
vin in 0 0v
vout out 0 0 


* NAND 

MP1 out_hp in vpmos vdd PMOS_32HP L=32n W=100n
MP2 out_hp in vpmos vdd PMOS_32HP L=32n W=100n
MN1 out_hp in dnmos 0 NMOS_32HP L=32n W=100n
MN2 dnmos in 0 0 NMOS_32HP L=32n W=100n


* Declarando o tipo de simulação 
.dc vin 0 2.5 0.01 vdd 0.5 2.5 0.5

*******************************************************************
* parametros de simulação

.control

run

* saida lógica
*spec 0 1K 100 3

    set color0=white
    set xbrushwidth=3

    plot v(out_hp) vs v(in)
    
.endc
.end