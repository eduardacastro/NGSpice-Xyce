*  cd ../../Users/Asus/Desktop/NGSpice/ckt-inversor/Xyce

.include "finfet.mod"

* Declaração das fontes
.param supply = 0.7
vdd vdd 0 dc 0.7

vin1 in1 0 PULSE (0 0. 0p 10p 10p 1200p 600p)
vin2 in2 0 PULSE (0 0. 0p 10p 10p 1200p 1200p)
vin3 in3 0 PULSE (0 0. 0p 10p 10p 1200p 600p)

Vagingp1 in1 inp1 dc -0.0445
Vagingp2 in2 inp2 dc -0.0397
Vagingp3 in3 inp3 dc -0.0397
Vagingn1 in1 inn1 dc 0.0445
Vagingn2 in2 inn2 dc 0.0425
Vagingn3 in3 inn3 dc 0.0445

.tran 0.001p 1000p
MP1 vpmos inp1 vdd vdd pmos_lvt L=20n NFIN=2 
MP2 out inp2 vpmos vpmos pmos_lvt L=20n NFIN=2
MP3 out inp3 vpmos vpmos pmos_lvt L=20n NFIN=2

MN1 out inn1 0 0 nmos_lvt L=20n NFIN=2
MN2 out inn2 v1nmos v1nmos nmos_lvt L=20n NFIN=2  
MN3 v1nmos inn3 0 0 nmos_lvt L=20n NFIN=2

*Variando In1
vaux out aux 0
* Positivo
*iexp 0 aux exp(0 34u 50p 2p 65p 4p)
* Negativo
iexp2 aux 0 exp(0 32u 50p 2p 65p 4p)


.OPTION OUTPUT INITIAL_INTERVAL=.1ps 350ps
.PRINT TRAN FORMAT=CSV v(out) v(in1) v(in2) v(in3)
.end