* Simulação de um inversor
* Incluindo o modelo do Transistor 
.include 32HP.mod
.include 32LP.mod

* Definindo a temperatura de operação
.TEMP 25


* Declarando parametros que serão utilizados nas simulações
.param supply = 0.9

* Declaração das fontes
valimentacao vdd 0 supply
vinput in 0 0.45
vout out 0 0
va 2 0 PULSE (0 1.8 0 0.1n 0.1n 10n 20n)
vb 2 0 PULSE (0 1.8 0 0.1n 0.1n 10n 20n)


MP1 vdd in1 out_32hp vdd pmos_32hp L=32n W=100n
MP2 vdd in2 out_32hp vdd pmos_32hp L=32n W=100n

MN1 out in1 mid_32hp vdd nmos_32hp L=32n W=100n
MN2 mid in2 gnd_32hp vdd nmos_32hp L=32n W=100n

* Declarando o tipo de simulação 
* .DC <fonte_que_sofrerá_variação> <valor_inicial_da_variação> <valor_final_da_variação> <passo_da_variação>
.dc vinput 0 0.9 0.01
*.dc vout 0 0.9 0.01 vinput 0 0.9 0.15

*******************************************************************
* parametros de simulação

.control

run

* saidas lógicas
plot out_32hp out_32lp


.endc