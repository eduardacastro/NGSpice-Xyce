*  cd ../../Users/Asus/Desktop/NGSpice/ckt-inversor/Xyce

.include "finfet.mod"
* Declaração das fontes
.param supply = 0.7
vdd vdd 0 dc 0.7
vin1 in2 0 PULSE (0 0.7 100p 10p 10p 1000p 1000p)
vin2 in1 0 PULSE (0 0.7 0p 10p 10p 300p 500p)
.tran 0.001p 1000p
Vagingp1 in1 inp1 dc -0.445
Vagingp2 in2 inp2 dc -0.445
Vagingn1 in1 inn1 dc 0.397
Vagingn2 in2 inn2 dc 0.445


MP1 out inp1 vdd vdd pmos_lvt L=20n NFIN=2 
MP2 out inp2 vdd vdd pmos_lvt L=20n NFIN=2
MN1 out inn1 dnmos 0 nmos_lvt L=20n NFIN=2 
MN2 dnmos inn2 0 0 nmos_lvt L=20n NFIN=2 




vaux out aux 0
* Positivo
iexp 0 aux exp(0 5u 200p 2p 215p 4p)
* Negativo
iexp2 aux 0 exp(0 5u 380p 2p 395p 4p)

.PRINT TRAN FORMAT=CSV v(out) v(in1) v(in2)
*Variando Inv1
.MEASURE TRAN HL TRIG v(in1) VAL='supply*0.5' RISE=2 TARG v(out) VAL='supply*0.5' FALL=2
.MEASURE TRAN LH TRIG v(in1) VAL='supply*0.5' FALL=1 TARG v(out) VAL='supply*0.5' RISE=1 
.MEASURE TRAN Fall TRIG v(out) VAL='supply*0.8' FALL=1 TARG v(out) VAL='supply*0.2' FALL=1
.MEASURE TRAN RISE TRIG v(out) VAL='supply*0.2' RISE=1 TARG v(out) VAL='supply*0.8' RISE=1

*Variando Inv2
*.MEASURE TRAN HL TRIG v(in2) VAL='supply*0.5' RISE=2 TARG v(out) VAL='supply*0.5' FALL=2
*.MEASURE TRAN LH TRIG v(in2) VAL='supply*0.5' FALL=1 TARG v(out) VAL='supply*0.5' RISE=1 
*.MEASURE TRAN Fall TRIG v(out) VAL='supply*0.8' FALL=1 TARG v(out) VAL='supply*0.2' FALL=1
*.MEASURE TRAN RISE TRIG v(out) VAL='supply*0.2' RISE=1 TARG v(out) VAL='supply*0.8' RISE=1

.end