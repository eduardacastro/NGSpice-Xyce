*  cd ../../NGSpice/ckt-inversor
* Definindo a temperatura de operação
.TEMP 25

.include "32HP.mod"

* Declaração das fontes
vdd vdd 0 dc 0.9
vin1 in 0 PULSE (0 0.9 100p 10p 10p 100p 300p)
.tran 0.001p 1000p


MP1 out in vdd vdd PMOS_32HP L=32n W=200n
MN1 out in 0 0 NMOS_32HP L=32n W=100n

.PRINT TRAN FORMAT=CSV v(out) v(in)
.MEASURE TRAN teste TRIG v(in) VAL=0.45 RISE=1 TARG v(out) VAL=0.45 FALL=1 

*meas tran tp_hl_in1 trig v(in1) val=0.45 rise=1 targ v(out) val=0.45 fall=1

.end