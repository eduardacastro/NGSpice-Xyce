*  cd ../../NGSpice/ckt-inversor
* Definindo a temperatura de operação
.TEMP 25

* Declarando parametros que serão utilizados nas simulações
.param agingp = -0.16
.param agingn = 0.16
.include 32HP.mod
* Declaração das fontes
vdd vdd 0 dc 0.9



vin1 in1 0 PULSE (0 0.9 100p 10p 10p 100p 300p)
Vagingp1 in1 inp1 dc -0.16
Vagingn1 in1 inn1 dc 0.16

MP1 out inp1 vdd vdd PMOS_32HP L=32n W=200n
MN1 out inn1 0 0 NMOS_32HP L=32n W=100n


*vaux out aux 0
* Positivo
*iexp 0 aux exp(0 145u 150p 2p 165p 4p)
* Negativo
*iexp2 aux 0 exp(0 155u 300p 2p 315p 4p)

*vaux out aux 0
*iexp 0 aux exp(0 200u 150p 2p 165p 4p)
*iexp2 aux 0 exp(0 190u 300p 2p 315p 4p)


.tran 0.001p 1000p
***********************
* parametros de simulação

.control
*  set color0=white
*  set xbrushwidth=3

*.plot v(outload2)-3 v(outload1)-2 v(outload)-1 v(out) v(in1)+1 

run
plot v(out) v(in1)+1
plot i(vdd)
meas tran tp_hl_in1 trig v(in1) val=0.45 rise=1 targ v(out) val=0.45 fall=1
meas tran tp_lh_in1 trig v(in1) val=0.45 fall=1 targ v(out) val=0.45 rise=1
meas tran tp_fall_in1 trig v(out) val=0.72 fall=1 targ v(out) val=0.18 fall=1
meas tran tp_rise_in1 trig v(out) val=0.18 rise=1 targ v(out) val=0.72 rise=1

.endc
.end