* Definindo a temperatura de operação
.TEMP 25

* Declarando parametros que serão utilizados nas simulações

.include 32LP.mod
.include 32HP.mod

* Declarando parametros que serão utilizados nas simulações
.param supply = 0.9

* Declaração das fontes
venable enable 0 0.45


* NAND 

MP1 out_nand enable vpmos vdd PMOS_32HP L=32n W=100n
MP2 out_nand out_oscilador vpmos vdd PMOS_32HP L=32n W=100n
MN1 out_nand enable dnmos 0 NMOS_32HP L=32n W=100n
MN2 dnmos out_oscilador 0 0 NMOS_32HP L=32n W=100n


* Declaração do inversor 1
MP_hp1 vdd out_nand out_inv1 vdd PMOS_32HP L=32n W=100n
MN_hp1 0   out_nand out_inv1 0   NMOS_32HP L=32n W=100n

* Declaração do inversor 2
MP_hp2 vdd out_inv1 out_inv2 vdd PMOS_32HP L=32n W=100n
MN_hp2 0   out_inv1 out_inv2 0   NMOS_32HP L=32n W=100n

* Declaração do inversor 3
MP_hp3 vdd out_inv2 out_inv3 vdd PMOS_32HP L=32n W=100n
MN_hp3 0   out_inv2 out_inv3 0   NMOS_32HP L=32n W=100n

* Declaração do inversor 4
MP_hp4 vdd out_inv2 out_inv4 vdd PMOS_32HP L=32n W=100n
MN_hp4 0   out_inv2 out_inv4 0   NMOS_32HP L=32n W=100n

* Declaração do inversor 5
MP_hp5 vdd out_inv4 out_inv5 vdd PMOS_32HP L=32n W=100n
MN_hp5 0   out_inv4 out_inv5 0   NMOS_32HP L=32n W=100n

* Declaração do inversor 6
MP_hp6 vdd out_inv5 out_inv6 vdd PMOS_32HP L=32n W=100n
MN_hp6 0   out_inv5 out_inv6 0   NMOS_32HP L=32n W=100n
* Declaração do inversor 7
MP_hp7 vdd out_inv6 out_inv7 vdd PMOS_32HP L=32n W=100n
MN_hp7 0   out_inv6 out_inv7 0   NMOS_32HP L=32n W=100n
* Declaração do inversor 8
MP_hp8 vdd out_inv7 out_inv8 vdd PMOS_32HP L=32n W=100n
MN_hp8 0   out_inv7 out_inv8 0   NMOS_32HP L=32n W=100n
* Declaração do inversor 9
MP_hp9 vdd out_inv8 out_inv9 vdd PMOS_32HP L=32n W=100n
MN_hp9 0   out_inv8 out_inv9 0   NMOS_32HP L=32n W=100n
* Declaração do inversor 10
MP_hp10 vdd out_inv9 out_inv10 vdd PMOS_32HP L=32n W=100n
MN_hp10 0   out_inv9 out_inv10 0   NMOS_32HP L=32n W=100n
* Declaração do inversor 11
MP_hp11 vdd out_inv10 out_oscilador vdd PMOS_32HP L=32n W=100n
MN_hp11 0   out_inv10 out_oscilador 0   NMOS_32HP L=32n W=100n


* Declarando o tipo de simulação 
.dc enable 0 0.9 0.01
*******************************************************************

.control

run

* saida lógica
*spec 0 1K 100 3

    set color0=white
    set xbrushwidth=3

    plot v(out_oscilador) 
    plot v(out_oscilador) v(enable)
    
.endc
.end