*  cd ../../NGSpice/ckt-nand
* Definindo a temperatura de operação
.TEMP 25

* Declarando parametros que serão utilizados nas simulações
.param agingp = -0.16
.param agingn = 0.16
.param Wp = 800n
.param Wn = 400n
.include 32HP.mod
* Declaração das fontes
vdd vdd 0 dc 0.9

* Variando Inv1
*vin1 in2 0 PULSE (0 0.9 300p 10p 10p 300p 600p)
*vin2 in1 0 PULSE (0 0.9 100p 10p 10p 2000p 4000p)


 
*Variando Inv2
vin1 in1 0 PULSE (0 0.9 100p 10p 10p 1000p 1000p)
vin2 in2 0 PULSE (0 0.9 0p 10p 10p 300p 500p)

Vagingp1 in1 inp1 dc agingp
Vagingn1 in1 inn1 dc agingn
Vagingp2 in2 inp2 dc agingp
Vagingn2 in2 inn2 dc agingn

MP1 out inp1 vdd vdd PMOS_32HP L=32n W=200n
MP2 out inp2 vdd vdd PMOS_32HP L=32n W=200n
MN1 out inn1 dnmos 0 NMOS_32HP L=32n W=100n
MN2 dnmos inn2 0 0 NMOS_32HP L=32n W=100n

*LOAD INV (FoF - Fanout of Four - emula 4 Invs usando sizing)
MPload outload out vdd vdd PMOS_32HP L=32n W=Wp
MNload outload out 0 0 NMOS_32HP L=32n W=Wn

MPloade1 outload1 outload vdd vdd PMOS_32HP L=32n W=Wp
MNloade1 outload1 outload 0 0 NMOS_32HP L=32n W=Wn

MPloade2 outload2 outload1 vdd vdd PMOS_32HP L=32n W=Wp
MNloade2 outload2 outload1 0 0 NMOS_32HP L=32n W=Wn

* variando in 1
vaux out aux 0
* sinal negativo
iexp aux 0 exp(0 160u 400p 2p 415p 4p)
*sinal positivo
iexp2 0 aux exp(0 105u 750p 2p 765p 4p)
* Declarando o tipo de simulação 

* variando in 2
*vaux out aux 0
* sinal negativo
*iexp aux 0 exp(0 150u 400p 2p 415p 4p)
*sinal positivo
*iexp2 0 aux exp(0 80u 650p 2p 665p 4p)
* Declarando o tipo de simulação 


*.tran 0.1p 500p
.tran 0.1p 900p
***********************
* parametros de simulação

.control

run
  set color0=gray
  set xbrushwidth=3
plot v(outload2)-3 v(outload1)-2 v(outload)-1 v(out) v(in1)+1 v(in2)+2 
*plot i(vaux)
*Variando Inv2
*meas tran tp_hl_in2_in1_0 trig v(in2) val=0.45 rise=1 targ v(out) val=0.45 fall=1
*meas tran tp_lh_in2_in1_0 trig v(in2) val=0.45 fall=1 targ v(out) val=0.45 rise=1
*meas tran tp_fall_in2_in1_0 trig v(out) val=0.72 fall=2 targ v(out) val=0.18 fall=2
*meas tran tp_rise_in2_in1_0 trig v(out) val=0.18 rise=2 targ v(out) val=0.72 rise=2

*Variando Inv1
meas tran tp_hl_in1_in2_0 trig v(in1) val=0.45 rise=2 targ v(out) val=0.45 fall=2
meas tran tp_lh_in1_in2_0 trig v(in1) val=0.45 fall=2 targ v(out) val=0.45 rise=2
meas tran tp_fall_in1_in2_0 trig v(out) val=0.72 fall=2 targ v(out) val=0.18 fall=2
meas tran tp_rise_in1_in2_0 trig v(out) val=0.18 rise=2 targ v(out) val=0.72 rise=2


.endc
.end