* Definindo a temperatura de operação
.TEMP 25

* Declarando parametros que serão utilizados nas simulações

.include 32HP.mod
* Declaração das fontes
vdd 1 0 dc 1.8

vin1 2 0 PULSE (0 1.8 0 0.1n 0.1n 5n 10n)
vin2 4 0 PULSE (0 1.8 0 0.1n 0.1n 10n 20n)

* Circuito da porta NAND
*<drain> <gate> <source> <bulk>
** portas em paralelo
*MP1 midsaida in1 vdd vdd PMOS_32HP L=32n W=100n
*MP2 midsaida in2 vdd vdd PMOS_32HP L=32n W=100n
MP1 3 2 1 1 PMOS_32HP L=32n W=100n
MP2 3 4 1 1 PMOS_32HP L=32n W=100n
MN1 3 2 5 0 NMOS_32HP L=32n W=100n
MN2 5 4 0 0 NMOS_32HP L=32n W=100n


** portas em série
*MN1 midsaida in1 mid mid NMOS_32HP L=32n W=100n
*MN2 mid in2 out out NMOS_32HP L=32n W=100n


* Declarando o tipo de simulação 
*.dc vin1 0 1.8 0.01
*.dc vin2 0 1.8 0.01 vin1 0 1.8 0.01
.tran 0.1n 50n
*******************************************************************
* parametros de simulação

.control

run

* saida lógica


.endc
.end