*  cd ../../Users/Asus/Desktop/NGSpice/ckt-inversor/Xyce
* Definindo a temperatura de operação
.include "finfet.mod"
.param supply = 0.7

* Declaração das fontes
vdd vdd 0 dc 0.7
vin1 in 0 PULSE (0 0.7 100p 10p 10p 300p 600p)
Vagingp1 in inp1 dc -0.445
Vagingn1 in inn1 dc 0.445
.tran 0.1p 1000p

 
MP1 out inp1 vdd vdd pmos_lvt L=20n NFIN=4
MN1 out inn1 0 0 nmos_lvt L=20n NFIN=4


vaux out aux 0
* Positivo
iexp 0 aux exp(0 10u 150p 2p 165p 4p)
* Negativo
vaux2 out aux2 0
iexp2 aux2 0 exp(0 5u 500p 2p 515p 4p)

.PRINT TRAN FORMAT=CSV v(out)
*.MEASURE TRAN HL TRIG v(in) VAL='supply*0.5' RISE=1 TARG v(out) VAL='supply*0.5' FALL=1 
*.MEASURE TRAN LH TRIG v(in) VAL='supply*0.5' FALL=1 TARG v(out) VAL='supply*0.5' RISE=1 
*.MEASURE TRAN Fall TRIG v(out) VAL='supply*0.8' FALL=1 TARG v(out) VAL='supply*0.2' FALL=1
*.MEASURE TRAN RISE TRIG v(out) VAL='supply*0.2' RISE=1 TARG v(out) VAL='supply*0.8' RISE=1

.end