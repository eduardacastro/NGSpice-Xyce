*  cd ../../Users/Asus/Desktop/NGSpice/ckt-oai/Xyce/oai-v1

.include "finfet.mod"

* Declaração das fontes
.param supply = 0.7
vdd vdd 0 dc 0.7
* Variando Inv1
vin1 in1 0 PULSE (0. 0. 0p 10p 10p 1200p 2400p)
vin2 in2 0 PULSE (0.7 0.7 0p 10p 10p 1200p 2400p)
vin3 in3 0 PULSE (0. 0. 0p 10p 10p 1200p 2400p)

.tran 0.001p 1000p

MP1 out in1 vdd vdd pmos_lvt L=20n NFIN=2
MP2 out in2 v1nmos v1nmos pmos_lvt L=20n NFIN=2  
MP3 v1nmos in3 vdd vdd pmos_lvt L=20n NFIN=2

MN1 out in1 vpmos vpmos nmos_lvt L=20n NFIN=2 
MN2 vpmos in2 0 0 nmos_lvt L=20n NFIN=2
MN3 vpmos in3 0 0 nmos_lvt L=20n NFIN=2

*Variando In1
vaux out aux 0
* Positivo
*iexp 0 aux exp(0 57u 350p 2p 365p 4p)
* Negativo
iexp2 aux 0 exp(0 49u 50p 2p 65p 4p)

.OPTION OUTPUT INITIAL_INTERVAL=.1ps 350ps
.PRINT TRAN FORMAT=CSV v(out) v(in1) v(in2) v(in3)
.end