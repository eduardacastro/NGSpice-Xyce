* Definindo a temperatura de operação
.TEMP 25

* Declarando parametros que serão utilizados nas simulações

.include 32LP.mod
.include 32HP.mod

* Declarando parametros que serão utilizados nas simulações
.param supply = 0.9

* Declaração das fontes
venable enable 0 PULSE (0 1.8 0 0.1n 0.1n 5n 10n)
vout_oscilador out_oscilador 0 PULSE (0 1.8 0 0.1n 0.1n 10n 20n)





* NAND 

MP1 out_nand enable vpmos vdd PMOS_32HP L=32n W=100n
MP2 out_nand out_oscilador vpmos vdd PMOS_32HP L=32n W=100n
MN1 out_nand enable dnmos 0 NMOS_32HP L=32n W=100n
MN2 dnmos out_oscilador 0 0 NMOS_32HP L=32n W=100n


* Declaração do inversor 1
MP_hp vdd out_nand out_inv1 vdd PMOS_32HP L=32n W=200n
MN_hp 0   out_nand out_inv1 0   NMOS_32HP L=32n W=100n

* Declaração do inversor 2
MP_hp vdd out_inv1 enable vdd PMOS_32HP L=32n W=200n
MN_hp 0   out_inv1 enable 0   NMOS_32HP L=32n W=100n

* Declarando o tipo de simulação 
.dc vinput 0 0.9 0.01
*******************************************************************
* parametros de simulação

.control

run

* saida lógica
*spec 0 1K 100 3

    set color0=white
    set xbrushwidth=3

    plot v(out_nand) v(out_lp) v(in)
    
.endc
.end