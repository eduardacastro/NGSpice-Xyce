* Definindo a temperatura de operação
.TEMP 25

* Declarando parametros que serão utilizados nas simulações
.param supply = 1.8
.include 32HP.mod
* Declaração das fontes
vdd vdd 0 supply
vout out 0 0
vmidsaida midsaida 0 0
vin1 2 0 PULSE (0 1.8 0 0.1n 0.1n 10n 20n)
vin2 2 0 PULSE (0 1.8 0 0.1n 0.1n 10n 20n)
* Modelagem dos transistores MOSFET
* PMOS com L=32nm e W=100nm
* NMOS com L=32nm e W=100nm



* Circuito da porta NAND
** portas em paralelo
MN1 vdd in1 midsaida  out NMOS_32HP L=32n W=100n
MN2 vdd in2 midsaida  out NMOS_32HP L=32n W=100n

** portas em série
MP1 midsaida in1 mid vdd PMOS_32HP L=32n W=100n
MP2 mid in2 0 vdd PMOS_32HP L=32n W=100n


* Declarando o tipo de simulação 
*.dc vin1 0 1.8 0.01
*.dc vin2 0 1.8 0.01 vin1 0 1.8 0.01
.tran 0.1n 100n
*******************************************************************
* parametros de simulação

.control

run

* saida lógica


.endc
.end