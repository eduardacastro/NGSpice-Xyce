* cd ../../NGSpice/ckt-oscilador_anel/cinco-portas
* Definindo a temperatura de operação
.TEMP 25

* Declarando parametros que serão utilizados nas simulações

.include 32LP.mod
.include 32HP.mod

* Declarando parametros que serão utilizados nas simulações
.param Wn = 100n
.param Wp = 200n
.param rad = 10u
* Declaração das fontes
vdd source 0 dc 0.9
venable enable 0 PWL(0 0 0.1n 0 0.11n 0.9) r=-1

.SUBCKT inv_32hp in out vdd gnd
iradp1 vdd out dc rad
iradn1 out gnd dc rad
MP_hp1 vdd in out vdd     PMOS_32HP L=32n W=Wp
MN_hp1 gnd in out gnd     NMOS_32HP L=32n W=Wn
.ends inv_32hp

.SUBCKT NAND A B out vdd gnd
iradp1 vdd out dc rad
iradp2 vdd out dc rad
iradn1 out dnmos dc rad
iradn2 dnmos gnd dc rad
*<drain gate source drain>
MP1 out A vdd vdd PMOS_32HP L=32n W=Wp
MP2 out B vdd vdd PMOS_32HP L=32n W=Wp
MN1 out A dnmos gnd NMOS_32HP L=32n W=Wn
MN2 dnmos B gnd gnd NMOS_32HP L=32n W=Wn
.ends NAND


* Xnand A B out vdd gnd NAND
Xnand enable out_oscilador out_nand source 0 NAND


* Xinv32hp in out vdd gnd inv_32hp
Xinv1 out_nand out_inv1 source 0 inv_32hp
Xinv2 out_inv1 out_inv2 source 0 inv_32hp
Xinv3 out_inv2 out_inv3 source 0 inv_32hp
Xinv4 out_inv3 out_inv4 source 0 inv_32hp
Xinv5 out_inv4 out_inv5 source 0 inv_32hp
Xinv6 out_inv5 out_inv6 source 0 inv_32hp
Xinv7 out_inv6 out_inv7 source 0 inv_32hp
Xinv8 out_inv7 out_inv8 source 0 inv_32hp
Xinv9 out_inv8 out_inv9 source 0 inv_32hp
Xinv10 out_inv9 out_inv10 source 0 inv_32hp
Xinv11 out_inv10 out_inv11 source 0 inv_32hp
Xinv12 out_inv11 out_inv12 source 0 inv_32hp
Xinv13 out_inv12 out_inv13 source 0 inv_32hp
Xinv14 out_inv13 out_inv14 source 0 inv_32hp
Xinv15 out_inv14 out_inv15 source 0 inv_32hp
Xinv16 out_inv15 out_oscilador source 0 inv_32hp


.tran 0.005n 2n
*******************************************************************

.control

run

* saida lógica
*spec 0 1K 100 3

    set color0=white
    set xbrushwidth=3

    *plot i(vaux)
    *plot v(out_inv2) 
    plot v(out_inv2) v(out_inv3)+1 v(out_inv4)+2 v(out_inv5)+3 v(out_inv1)+4 
    
    *plot v(out_inv2) v(out_inv1)
    MEAS TRAN periodo TRIG v(out_inv2) VAL=0.45 RISE=2 TARG v(out_inv2) VAL=0.45 RISE=3
    MEAS TRAN tempo_alto TRIG v(out_inv2) VAL=0.45 RISE=2 TARG v(out_inv2) VAL=0.45 FALL=3
    MEAS TRAN tempo_baixo TRIG v(out_inv2) VAL=0.45 FALL=3 TARG v(out_inv2) VAL=0.45 RISE=3
    MEAS TRAN trise TRIG v(out_inv2) VAL=0.18 RISE=2 TARG v(out_inv2) VAL=0.72 RISE=2
    MEAS TRAN tfall TRIG v(out_inv2) VAL=0.72 FALL=2 TARG v(out_inv2) VAL=0.18 FALL=2
.endc
.end