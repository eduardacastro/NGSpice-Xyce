*  cd ../../Users/Asus/Desktop/NGSpice/ckt-inversor/Xyce
* Definindo a temperatura de operação
.include "finfet.mod"
.param supply = 0.7

* Declaração das fontes
vdd vdd 0 dc 0.7
vin1 in 0 PULSE (0.7 0.7 0p 10p 10p 100p 2400p)
.tran 0.001p 1000p

 
MP1 out in vdd vdd pmos_lvt L=20n NFIN=2
MN1 out in 0 0 nmos_lvt L=20n NFIN=2


*  SET
************
vaux out aux 0
* Positivo
iexp 0 aux exp(0 63u 50p 2p 65p 4p)
* Negativo
*iexp2 aux 0 exp(0 50u 550p 2p 565p 4p)



.OPTION OUTPUT INITIAL_INTERVAL=.1ps 350ps
.PRINT TRAN FORMAT=CSV v(out) v(in)

.end