*  cd ../../Users/Asus/Desktop/NGSpice/ckt-inversor
* Definindo a temperatura de operação
.TEMP 25
.param agingp = -0.16
.param agingn = 0.16
.include "32HP.mod"

* Declaração das fontes
vdd vdd 0 dc 0.9
vin1 in 0 PULSE (0 0.9 100p 10p 10p 100p 300p)
Vagingp1 inp1 in dc 0.16
Vagingn1 in inn1 dc 0.16
.tran 0.001p 1000p


MP1 out inp1 vdd vdd PMOS_32HP L=32n W=200n
MN1 out inn1 0 0 NMOS_32HP L=32n W=100n

vaux out aux 0
* Positivo
iexp 0 aux exp(0 145u 150p 2p 165p 4p)
* Negativo
iexp2 aux 0 exp(0 155u 300p 2p 315p 4p)

.PRINT TRAN FORMAT=CSV v(out) v(in)
.MEASURE TRAN HL TRIG v(in) VAL=0.45 RISE=1 TARG v(out) VAL=0.45 FALL=1 
.MEASURE TRAN LH TRIG v(in) VAL=0.45 FALL=1 TARG v(out) VAL=0.45 RISE=1 
.MEASURE TRAN Fall TRIG v(out) VAL=0.72 FALL=1 TARG v(out) VAL=0.18 FALL=1
.MEASURE TRAN RISE TRIG v(out) VAL=0.18 RISE=1 TARG v(out) VAL=0.72 RISE=1

*meas tran tp_hl_in1 trig v(in1) val=0.45 rise=1 targ v(out) val=0.45 fall=1
*meas tran tp_lh_in1 trig v(in1) val=0.45 fall=1 targ v(out) val=0.45 rise=1
*meas tran tp_fall_in1 trig v(out) val=0.72 fall=1 targ v(out) val=0.18 fall=1
*meas tran tp_rise_in1 trig v(out) val=0.18 rise=1 targ v(out) val=0.72 rise=1

.end