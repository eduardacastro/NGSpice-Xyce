* Definindo a temperatura de operação
.TEMP 25

* Declarando parametros que serão utilizados nas simulações

.include 32HP.mod
* Declaração das fontes
vdd vdd 0 dc 0.9

*vin1 in1 0 PULSE (0 0.9 0 0.1n 0.1n 5n 10n)
*vin2 in2 0 PULSE (0 0.9 0 0.1n 0.1n 10n 20n)

vin1 in1 0 PULSE (0 0.9 300p 10p 10p 100p 10n)
vin2 in2 0 PULSE (0 0.9 100p 10p 10p 100p 20n)



MP1 out in1 vpmos vdd PMOS_32HP L=32n W=100n
MP2 out in2 vpmos vdd PMOS_32HP L=32n W=100n
MN1 out in1 dnmos 0 NMOS_32HP L=32n W=100n
MN2 dnmos in2 0 0 NMOS_32HP L=32n W=100n


.tran 0.1p 500p
***********************
* parametros de simulação

.control

run
plot v(out) v(in1)+1 v(in2)
meas tran tp_hl_in2_in1_0 trig v(in2) val=0.45 rise=1 targ v(out) val=0.45 fall=1
meas tran tp_lh_in2_in1_0 trig v(in2) val=0.45 fall=1 targ v(out) val=0.45 rise=1
meas tran tp_hl_in1_in2_0 trig v(in1) val=0.45 rise=1 targ v(out) val=0.45 fall=2
meas tran tp_lh_in1_in2_0 trig v(in1) val=0.45 fall=1 targ v(out) val=0.45 rise=2
meas tran tp_fall_in2_in1_0 trig v(out) val=0.72 fall=1 targ v(out) val=0.18 fall=1
meas tran tp_rise_in2_in1_0 trig v(out) val=0.18 rise=1 targ v(out) val=0.72 rise=1
meas tran tp_fall_in2_in1_0 trig v(out) val=0.72 fall=2 targ v(out) val=0.18 fall=2
meas tran tp_rise_in2_in1_0 trig v(out) val=0.18 rise=2 targ v(out) val=0.72 rise=2

.endc
.end