*  cd ../../Users/Asus/Desktop/NGSpice/ckt-inversor/Xyce
* Definindo a temperatura de operação
.include "finfet.mod"
.param supply = 0.7

* Declaração das fontes
vdd vdd 0 dc 0.7
vin1 in 0 PULSE (0 0.7 100p 10p 10p 100p 300p)
.tran 0.001p 1000p

 
MP1 out in vdd vdd pmos_lvt L=20n W=54n NFIN=4
MN1 out in 0 0 nmos_lvt L=20n W=54n NFIN=4

*cload out 0 0.5f

.PRINT TRAN FORMAT=CSV v(out) v(in)
.MEASURE TRAN HL TRIG v(in) VAL='supply*0.5' RISE=1 TARG v(out) VAL='supply*0.5' FALL=1 
.MEASURE TRAN LH TRIG v(in) VAL='supply*0.5' FALL=1 TARG v(out) VAL='supply*0.5' RISE=1 
.MEASURE TRAN Fall TRIG v(out) VAL='supply*0.8' FALL=1 TARG v(out) VAL='supply*0.2' FALL=1
.MEASURE TRAN RISE TRIG v(out) VAL='supply*0.2' RISE=1 TARG v(out) VAL='supply*0.8' RISE=1

.end