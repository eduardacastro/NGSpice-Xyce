Simulação_transiente_de_um_Inversor
*
* Detalher sobre o Ckt
*
* Copyright (c) 2023 - Eduarda de Castro Guterres
* Distribuição sob a licença GNU GPLv2 
*
****************************************************************
*Incluindo os modelos de transistores
.include 32_HP.mod
.include 32_LP.mod

* Def. da Temperatura
.TEMP 25

****************************************************************
*Parametro que será utilizado na simulação
.param supply = 0.9

* Descrição das fontes
vSignal vdd  0  0.9
vinput  in   0  PULSE( 0 0.9 1n 1p 1p 1n 2n) 

* Inversor
MP vdd in out vdd PMOS_hp L=32n W=100n
MN 0   in out 0   NMOS_hp L=32n W=100n

* Capacitancia de saída para emular uma carga
Cload out 0 5f

****************************************************************
* Parametros da Simulação

.tran 0.1p 32n

*Comandos measure para a realização de medidas
.MEAS TRAN integral_vdd INTEG v(vSignal) from=0.9n to 1.1n
.MEAS TRAN integral_in  INTEG v(vinput) from=0.9n to 1.1n

.MEAS TRAN tp_lh   TRIG v(in)  val=0.5 FALL=1 TARG v(out) val=0.5 RISE=1
.MEAS TRAN tp_hl   TRIG v(in)  val=0.5 RISE=1 TARG v(out) val=0.5 FALL=1
.MEAS TRAN tp_fall TRIG v(out) val=0.75 FALL=1 TARG v(out) val=0.25 FALL=1
.MEAS TRAN tp_rise TRIG v(out) val=0.25 RISE=1 TARG v(out) val=0.75 RISE=1