Simulacao_transiente_de_um_Inversor
*
* Detalher sobre o Ckt
*
* Copyright (c) 2023 - Eduarda de Castro Guterres
* Distribuicao sob a licenca GNU GPLv2 
*
****************************************************************
*Incluindo os modelos de transistores
.include 32HP.mod
.include 32LP.mod

* Def. da Temperatura
.TEMP 25

****************************************************************
*Parametro que sera utilizado na simulacao
.param supply = 0.9

* Descricao das fontes
valimentacao vdd 0 0.9
vinput in 0 PULSE (0 0.9 1n 1p 1p 1n 2n) 

* Inversor
MP vdd in out vdd PMOS_32hp L=32n W=100n
MN 0 in out 0 NMOS_32hp L=32n W=100n

* Capacitancia de saida para emular uma carga
Cload out 0 5f

****************************************************************
* Parametros da Simulacao

.tran 0.1p 3n

*Comandos measure para a realizacao de medidas
*.MEAS TRAN integral_vdd INTEG i(valimentacao) from=1.9n to=2.2n
.MEAS TRAN integral_in1 INTEG i(vinput) from=0.9n to=1.1n
.MEAS TRAN integral_in2 INTEG i(vinput) from=1.9n to=2.1n

*.MEAS TRAN tp_lh TRIG v(in) val=0.5 FALL=1 TARG v(out) val=0.5 RISE=1
*.MEAS TRAN tp_hl TRIG v(in) val=0.5 RISE=1 TARG v(out) val=0.5 FALL=1
*.MEAS TRAN tp_fall TRIG v(out) val=0.75 FALL=1 TARG v(out) val=0.25 FALL=1
*.MEAS TRAN tp_rise TRIG v(out) val=0.25 RISE=1 TARG v(out) val=0.75 RISE=1

.end