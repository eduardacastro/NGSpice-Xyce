*  cd ../../NGSpice/ckt-inversor
* Definindo a temperatura de operação
.TEMP 25

* Declarando parametros que serão utilizados nas simulações
.param agingp = -0.16
.param agingn = 0.16
.include 32HP.mod
* Declaração das fontes
vdd vdd 0 dc 0.9



vin1 in1 0 PULSE (0 0.9 100p 10p 10p 100p 300p)
Vagingp1 in1 inp1 dc agingp
Vagingn1 in1 inn1 dc agingn

MP1 out inp1 vdd vdd PMOS_32HP L=32n W=200n
MN1 out inn1 0 0 NMOS_32HP L=32n W=100n


*LOAD INV (FoF - Fanout of Four - emula 4 Invs usando sizing)
MPload outload out vdd vdd PMOS_32HP L=32n W=800n
MNload outload out 0 0 NMOS_32HP L=32n W=400n

MPloade1 outload1 outload vdd vdd PMOS_32HP L=32n W=800n
MNloade1 outload1 outload 0 0 NMOS_32HP L=32n W=400n

MPloade2 outload2 outload1 vdd vdd PMOS_32HP L=32n W=800n
MNloade2 outload2 outload1 0 0 NMOS_32HP L=32n W=400n

vaux out aux 0
iexp 0 aux exp(0 140u 150p 2p 165p 4p)
iexp2 aux 0 exp(0 150u 300p 2p 315p 4p)

*vaux out aux 0
*iexp 0 aux exp(0 200u 150p 2p 165p 4p)
*iexp2 aux 0 exp(0 190u 300p 2p 315p 4p)


.tran 0.1p 600p
***********************
* parametros de simulação

.control
  set color0=white
  set xbrushwidth=3

  plot v(outload2)-3 v(outload1)-2 v(outload)-1 v(out) v(in1)+1 

run
*plot v(out) v(in1)+1
*plot i(vdd)
meas tran tp_hl_in1 trig v(in1) val=0.45 rise=1 targ v(out) val=0.45 fall=1
meas tran tp_lh_in1 trig v(in1) val=0.45 fall=1 targ v(out) val=0.45 rise=1
meas tran tp_fall_in1 trig v(out) val=0.72 fall=1 targ v(out) val=0.18 fall=1
meas tran tp_rise_in1 trig v(out) val=0.18 rise=1 targ v(out) val=0.72 rise=1

.endc
.end