*  cd ../../Users/Asus/Desktop/NGSpice/ckt-inversor/Xyce

.include "finfet.mod"

* Declaração das fontes
.param supply = 0.7
vdd vdd 0 dc 0.7
vin2 in4 0 PULSE (0 0.7 0p 10p 10p 300p 500p)
vin1 in2 0 PULSE (0 0.7 100p 10p 10p 1000p 1000p)
vin3 in1 0 PULSE (0 0.7 100p 10p 10p 1000p 1000p)
vin4 in3 0 PULSE (0 0.7 100p 10p 10p 1000p 1000p)

.tran 0.001p 1000p


MP1 out in1 vdd vdd pmos_lvt L=20n NFIN=2 
MP2 out in2 vdd vdd pmos_lvt L=20n NFIN=2
MP3 out in3 vdd vdd pmos_lvt L=20n NFIN=2
MP4 out in4 vdd vdd pmos_lvt L=20n NFIN=2

MN1 out in1 v2nmos v2nmos nmos_lvt L=20n NFIN=2
MN2 v2nmos in2 v3nmos v3nmos nmos_lvt L=20n NFIN=2  
MN3 v3nmos in3  v4nmos v4nmos nmos_lvt L=20n NFIN=2 
MN4 v4nmos in4 0 0 nmos_lvt L=20n NFIN=2 


.OPTION OUTPUT INITIAL_INTERVAL=.1ps 350ps
.PRINT TRAN FORMAT=CSV v(out) v(in1) v(in2) v(in3)

*Variando Inv1
.MEASURE TRAN HL1 TRIG v(in1) VAL='supply*0.5' RISE=2 TARG v(out) VAL='supply*0.5' FALL=2
.MEASURE TRAN LH1 TRIG v(in1) VAL='supply*0.5' FALL=1 TARG v(out) VAL='supply*0.5' RISE=1

*Variando Inv2
.MEASURE TRAN HL2 TRIG v(in2) VAL='supply*0.5' RISE=2 TARG v(out) VAL='supply*0.5' FALL=2
.MEASURE TRAN LH2 TRIG v(in2) VAL='supply*0.5' FALL=1 TARG v(out) VAL='supply*0.5' RISE=1

*Variando Inv3
.MEASURE TRAN HL3 TRIG v(in3) VAL='supply*0.5' RISE=2 TARG v(out) VAL='supply*0.5' FALL=2
.MEASURE TRAN LH3 TRIG v(in3) VAL='supply*0.5' FALL=1 TARG v(out) VAL='supply*0.5' RISE=1

*Variando Inv3
.MEASURE TRAN HL4 TRIG v(in4) VAL='supply*0.5' RISE=2 TARG v(out) VAL='supply*0.5' FALL=2
.MEASURE TRAN LH4 TRIG v(in4) VAL='supply*0.5' FALL=1 TARG v(out) VAL='supply*0.5' RISE=1


.MEASURE TRAN Fall2 TRIG v(out) VAL='supply*0.8' FALL=2 TARG v(out) VAL='supply*0.2' FALL=2
.MEASURE TRAN RISE2 TRIG v(out) VAL='supply*0.2' RISE=2 TARG v(out) VAL='supply*0.8' RISE=2

.end