* Definindo a temperatura de operação
.TEMP 25

* Declarando parametros que serão utilizados nas simulações

.include 32LP.mod
.include 32HP.mod

* Declarando parametros que serão utilizados nas simulações
.param supply = 0.9

* Declaração das fontes
vdd source 0 dc 0.9
venable enable 0 PWL(0 0.9) r=-1
*vclock 7 5 PWL(0 1 20ns 0) r=-1

* NAND 
MP1 out_nand enable        source   source PMOS_32HP L=32n W=100n
MP2 out_nand out_oscilador source   source PMOS_32HP L=32n W=100n
MN1 out_nand enable        dnmos    0      NMOS_32HP L=32n W=100n
MN2 dnmos    out_oscilador 0        0      NMOS_32HP L=32n W=100n  


.SUBCKT inv_32hp in out vdd gnd
MP_hp1 vdd in out vdd     PMOS_32HP L=32n W=100n
MN_hp1 gnd in out gnd     NMOS_32HP L=32n W=100n
.ends inv_32hp

* Xinv32hp in out vdd gnd inv_32hp
Xinv1 out_oscilador out_inv1 source 0 inv_32hp
X2inv2 out_inv1 out_oscilador source 0 inv_32hp



* Declarando o tipo de simulação 

.tran 0.005n 1n
*******************************************************************

.control

run

* saida lógica
*spec 0 1K 100 3

    set color0=white
    set xbrushwidth=3

    plot v(out_oscilador) 
    plot v(out_oscilador) v(enable)
    
.endc
.end