* Simulação de um inversor
* Incluindo o modelo do Transistor 
.include 32HP.mod
.include 32LP.mod

* Definindo a temperatura de operação
.TEMP 25

* Declarando parametros que serão utilizados nas simulações
.param supply = 0.9

* Declaração das fontes
valimentacao vdd 0 supply
vinput in 0 0.45
vout out 0 0

vpmos_b dpmos_b out 0
vnmos_b out dnmos_b 0

vpmos_a out dpmos_a 0
vnmos_a out dnmos_a 0

* Declaração do inversor
MP vdd in out_32hp vdd pmos_32hp L=32n W=200n
MN 0   in out_32hp 0   nmos_32hp L=32n W=100n

MP_lp vdd in out_32lp vdd PMOS_32lp L=32n W=200n
MN_lp 0   in out_32lp 0   NMOS_32lp L=32n W=100n

* Pb vdd in dpmos_b vdd PMOS_1p L=32n W=200n
* MNb 0   in dnmos_b 0   NMOS_1p L=32n W=100n

* Pa vdd in dpmos_a vdd PMOS_1p L=32n W=200n
* MNa 0   in dnmos_a 0   NMOS_1p L=32n W=100n

* Declarando o tipo de simulação 
* .DC <fonte_que_sofrerá_variação> <valor_inicial_da_variação> <valor_final_da_variação> <passo_da_variação>
.dc vinput 0 0.9 0.01
*dc vout 0 0.9 -/01 vinput 0 0.9 0.15

.end