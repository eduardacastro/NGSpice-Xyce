*  cd ../../Users/Asus/Desktop/NGSpice/ckt-nor/Xyce/nor-2

.include "finfet.mod"
.param supply = 0.7
* Declaração das fontes
vdd vdd 0 dc 0.7
vin1 in2 0 PULSE (0 0.0 100p 10p 10p 1000p 1000p)
vin2 in1 0 PULSE (0 0.7 0p 10p 10p 300p 500p)
.tran 0.001p 1000p
Vagingp1 in1 inp1 dc -0.0445
Vagingp2 in2 inp2 dc -0.0397
Vagingn1 in1 inn1 dc 0.0445
Vagingn2 in2 inn2 dc 0.0445



MP1 out inp1 vpmos vdd pmos_lvt L=20n NFIN=2 
MP2 vpmos inp2 vdd vdd pmos_lvt L=20n NFIN=2 
MN1 out inn1 0 0 nmos_lvt L=20n NFIN=2 
MN2 out inn2 0 0 nmos_lvt L=20n NFIN=2 

vaux out aux 0
* Positivo
iexp 0 aux exp(0 60u 150p 2p 165p 4p)
* Negativo
iexp2 aux 0 exp(0 25u 350p 2p 365p 4p)

.OPTION OUTPUT INITIAL_INTERVAL=.1ps 350ps
.PRINT TRAN FORMAT=CSV v(out) v(in1) v(in2)

.end