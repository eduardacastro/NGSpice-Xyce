* cd ../../NGSpice/ckt-oscilador_anel/treze-porta
* Definindo a temperatura de operação
.TEMP 25

* Declarando parametros que serão utilizados nas simulações

.include 32LP.mod
.include 32HP.mod

* Declarando parametros que serão utilizados nas simulações
.param Wn = 100n
.param Wp = 200n


* Declaração das fontes
vdd source 0 dc 0.9
venable enable 0 PWL(0 0 0.1n 0 0.11n 0.9) r=-1
*vclock 7 5 PWL(0 1 20ns 0) r=-1

.SUBCKT inv_32hp in out vdd gnd
iradp1 vdd out dc -10000n
iradn1 gnd out dc 10000n

MP_hp1 vdd in out vdd     PMOS_32HP L=32n W=Wp
MN_hp1 gnd in out gnd     NMOS_32HP L=32n W=Wn
.ends inv_32hp

.SUBCKT NAND A B out vdd gnd
iradp1 vdd out dc -10000n
iradp2 vdd out dc -10000n
iradn1 dnmos out dc 10000n
iradn2 gnd dnmos dc 10000n
*<drain gate source drain>
MP1 out A vdd vdd PMOS_32HP L=32n W=150n
MP2 out B vdd vdd PMOS_32HP L=32n W=150n
MN1 out A dnmos gnd NMOS_32HP L=32n W=250n
MN2 dnmos B gnd gnd NMOS_32HP L=32n W=250n
.ends NAND

* Xnand A B out vdd gnd NAND
Xnand enable out_oscilador out_nand source 0 NAND


* Xinv32hp in out vdd gnd inv_32hp
Xinv1 out_nand out_inv1 source 0 inv_32hp
Xinv2 out_inv1 out_inv2 source 0 inv_32hp
Xinv3 out_inv2 out_inv3 source 0 inv_32hp
Xinv4 out_inv3 out_inv4 source 0 inv_32hp
Xinv5 out_inv4 out_inv5 source 0 inv_32hp
Xinv6 out_inv5 out_inv6 source 0 inv_32hp
Xinv7 out_inv6 out_inv7 source 0 inv_32hp
Xinv8 out_inv7 out_inv8 source 0 inv_32hp
Xinv9 out_inv8 out_inv9 source 0 inv_32hp
Xinv10 out_inv9 out_inv10 source 0 inv_32hp
Xinv11 out_inv10 out_inv11 source 0 inv_32hp
Xinv12 out_inv11 out_oscilador source 0 inv_32hp

****************************************************************************
* Saida do Oscilador
* Declaração do inversor 5
*MP_hp17 out_inv17 out_oscilador source source PMOS_32HP L=32n W=80n
*MN_hp17 out_inv17 out_oscilador 0      0      NMOS_32HP L=32n W=100n

* Declaração do inversor 5
*MP_hp18 out_inv18 out_inv17 source source PMOS_32HP L=32n W=200n
*MN_hp18 out_inv18 out_inv17 0      0      NMOS_32HP L=32n W=100n

* Declaração do inversor 5
*MP_hp19 out_inv19 out_inv18 source source PMOS_32HP L=32n W=150n
*MN_hp19 out_inv19 out_inv18 0      0      NMOS_32HP L=32n W=8000n



* Declarando o tipo de simulação 

.tran 0.005n 1n
*******************************************************************

.control

run

* saida lógica
*spec 0 1K 100 3

    set color0=white
    set xbrushwidth=3

    plot v(out_inv2) 
    plot v(out_inv2) v(enable)
    MEAS TRAN periodo TRIG v(out_inv2) VAL=0.45 RISE=2 TARG v(out_inv2) VAL=0.45 RISE=3
    MEAS TRAN tempo_alto TRIG v(out_inv2) VAL=0.45 RISE=2 TARG v(out_inv2) VAL=0.45 FALL=3
    MEAS TRAN tempo_baixo TRIG v(out_inv2) VAL=0.45 FALL=3 TARG v(out_inv2) VAL=0.45 RISE=3
    MEAS TRAN trise TRIG v(out_inv2) VAL=0.18 RISE=2 TARG v(out_inv2) VAL=0.72 RISE=2
    MEAS TRAN tfall TRIG v(out_inv2) VAL=0.72 FALL=2 TARG v(out_inv2) VAL=0.18 FALL=2
.endc
.end