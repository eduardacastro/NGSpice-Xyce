* cd ../../NGSpice/ckt-nand
* Definindo a temperatura de operação
.TEMP 25

* Declarando parametros que serão utilizados nas simulações

.include 32HP.mod
* Declaração das fontes
vdd vdd 0 dc 1.8

vin1 in1 0 PULSE (0 1.8 0 0.1n 0.1n 5n 10n)
vin2 in2 0 PULSE (0 1.8 0 0.1n 0.1n 10n 20n)

; Adicione uma fonte de tensão após in1
vfontep1 in1 vfontep1 dc -0.16
vfontep2 in2 vfontep2 dc -0.16
vfonten1 in1 vfonten1 dc 0.16
vfonten2 in2 vfonten2 dc 0.16
* Circuito da porta NAND
*<drain> <gate> <source> <bulk>
** portas em paralelo
*MP1 midsaida in1 vdd vdd PMOS_32HP L=32n W=100n
*MP2 midsaida in2 vdd vdd PMOS_32HP L=32n W=100n
MP1 out vfontep1 vdd vdd PMOS_32HP L=32n W=100n
MP2 out vfontep2 vdd vdd PMOS_32HP L=32n W=100n
MN1 out vfonten1 dnmos 0 NMOS_32HP L=32n W=100n
MN2 dnmos vfonten2 0 0 NMOS_32HP L=32n W=100n


** portas em série
*MN1 midsaida in1 mid mid NMOS_32HP L=32n W=100n
*MN2 mid in2 out out NMOS_32HP L=32n W=100n


* Declarando o tipo de simulação 
*.dc vin1 0 1.8 0.01
*.dc vin2 0 1.8 0.01 vin1 0 1.8 0.01
.tran 1n 50n
***********************
* parametros de simulação

.control

run
 set color0=white
    set xbrushwidth=3
* saida lógica
spec 0 1K 100 3
*plot v(out) v(in1) v(in2)
plot v(in1) v(in2)
plot v(out)
fft v(out)
plot mag(v(out))

.endc
.end